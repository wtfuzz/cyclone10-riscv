@00000000
91000537
00050513
0FF00293
00550223
00550A23
00300293
00550023
900005B7
00058593
08300293
005581A3
00000293
005580A3
01B00293
00558023
00300293
005581A3
04100393
00758023
00100337
00000E13
01C50023
001E0E13
04100393
00758023
000073B3
00138393
FE731EE3
FE5FF06F
	 
