@00000000
37 06 00 91 13 06 06 00 93 02 F0 0F 23 02 56 00
23 0A 56 00 93 02 10 00 23 00 56 00 6F F0 5F FE
13 01 00 0D E7 00 01 00 13 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
23 2E 11 FE 23 2C 51 FE 23 2A 61 FE 23 28 71 FE
23 26 A1 FE 23 24 B1 FE 23 22 C1 FE 23 20 D1 FE
23 2E E1 FC 23 2C F1 FC 23 2A 01 FD 23 28 11 FD
23 26 C1 FD 23 24 D1 FD 23 22 E1 FD 23 20 F1 FD
13 01 01 FC EF 00 00 5D 83 20 C1 03 83 22 81 03
03 23 41 03 83 23 01 03 03 25 C1 02 83 25 81 02
03 26 41 02 83 26 01 02 03 27 C1 01 83 27 81 01
03 28 41 01 83 28 01 01 03 2E C1 00 83 2E 81 00
03 2F 41 00 83 2F 01 00 13 01 01 04 73 00 20 30
97 11 00 00 93 81 01 D6 13 01 00 63 37 06 00 91
13 06 06 00 93 02 20 00 23 00 56 00 13 05 80 63
93 05 80 63 63 08 B5 00 23 20 05 00 13 05 45 00
6F F0 5F FF 93 02 30 00 23 00 56 00 13 05 C0 65
13 01 C1 FF 93 05 C0 65 63 0E B5 00 83 26 05 00
13 05 45 00 23 20 A1 00 E7 80 06 00 03 25 01 00
6F F0 5F FE 93 02 40 00 23 00 56 00 13 01 41 00
93 02 50 00 23 00 56 00 B7 05 00 90 93 85 05 00
93 02 30 08 A3 81 55 00 93 02 00 00 A3 80 55 00
93 02 B0 01 23 80 55 00 93 02 30 00 A3 81 55 00
93 03 E0 02 23 80 75 00 EF 00 40 09 6F 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 6F 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00
@00000630
00 00 00 90 00 00 00 91
@00000638
83 47 05 00 63 94 07 00 67 80 00 00 83 26 00 63
13 05 15 00 23 80 F6 00 6F F0 9F FE 67 80 00 00
@00000658
6F 00 00 00
