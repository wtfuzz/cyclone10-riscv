@00000000
91000637
00060613
0FF00293
00560223
00560A23
00100293
00560023
0D000113
000100E7
00000013
00000000
00000000
00000000
00000000
00000000
00000000
FE112E23
FE512C23
FE612A23
FE712823
FEA12623
FEB12423
FEC12223
FED12023
FCE12E23
FCF12C23
FD012A23
FD112823
FDC12623
FDD12423
FDE12223
FDF12023
FC010113
180000EF
03C12083
03812283
03412303
03012383
02C12503
02812583
02412603
02012683
01C12703
01812783
01412803
01012883
00C12E03
00812E83
00412F03
00012F83
04010113
30200073
00002197
1C018193
80000117
12810113
91000637
00060613
00200293
00560023
80000517
11050513
80000597
11058593
00B50863
00052023
00450513
FF5FF06F
00300293
00560023
80000517
0F050513
FFC10113
80000597
0E458593
00B50E63
00052683
00450513
00A12023
000680E7
00012503
FE1FF06F
00400293
00560023
00410113
00500293
00560023
900005B7
00058593
08300293
005581A3
00000293
005580A3
01B00293
00558023
00300293
005581A3
02E00393
00758023
544010EF
0000006F
00000000
00000000
FE010113
00812E23
02010413
FEA42623
FEC42703
000017B7
38878793
02F707B3
FEF42623
0100006F
FEC42783
FFF78793
FEF42623
FEC42783
FE0798E3
00000013
00000013
01C12403
02010113
00008067
90000737
00574783
0407F793
FE078CE3
00B70023
00008067
00008067
FC010113
03512223
03612023
00C62A83
01062B03
02812C23
02912A23
03212823
03312623
03412423
01712E23
02112E23
01812C23
01912A23
01A12823
01B12623
00050913
00058993
00060A13
00000B93
00100493
00000413
00048613
00040693
00090513
00098593
0C1000EF
04BB9C63
05557A63
00000B93
00900C93
0084E7B3
04079C63
000B0023
03C12083
03812403
03412483
03012903
02C12983
02812A03
02412A83
02012B03
01C12B83
01812C03
01412C83
01012D03
00C12D83
04010113
00008067
035407B3
0354B433
035484B3
00878433
F85FF06F
00048613
00040693
00090513
00098593
041000EF
00048613
00040693
00098593
00050A93
00050D13
00090513
5FD000EF
00CA2C03
00050913
00058993
000C0613
00000693
00048513
00040593
005000EF
000B9E63
01504C63
00041463
0584E063
00050493
00058413
F3DFF06F
03000793
01ACDC63
000A4703
03700793
00477713
00071463
05700793
015787B3
00FB0023
001B8B93
001B0B13
FC9FF06F
03000793
FE9FF06F
0105A703
00C5A683
00100793
02F55633
00D67C63
00000693
00900893
00079A63
00070023
00008067
02D787B3
FE1FF06F
00C5A803
02F55633
0307D333
02F57533
00069A63
00C04863
0307EE63
00030793
FCDFF06F
03000793
00C8DC63
0005C803
03700793
00487813
00081463
05700793
00C787B3
00F70023
00168693
00170713
FCDFF06F
03000793
FE9FF06F
FE010113
00812C23
01062783
00462403
00912A23
01312623
01412423
00112E23
01212823
00050993
00058A13
00060493
0007C703
00178793
00070463
0E804063
0084C783
00078463
FFF40413
0004C783
0027F793
00078A63
00C4A783
01000713
0CE79263
FFE40413
0004A783
00040913
0097F793
0C078863
0084C583
00058663
00098513
000A00E7
0004C783
0027F793
02078C63
00C4A783
01000713
0CE79063
03000593
00098513
000A00E7
0004C783
05800593
0047F793
00079463
07800593
00098513
000A00E7
0004C783
00040913
0017F793
0A079463
0104A903
00094583
00190913
0A059863
0004A783
00800713
0097F793
00E79463
0A804463
01C12083
01812403
01412483
01012903
00C12983
00812A03
02010113
00008067
FFF40413
F11FF06F
00800713
F4E790E3
FFF40413
F39FF06F
02000593
00098513
000A00E7
FFF90913
FF2048E3
FFF40793
00045463
00000413
40878433
F21FF06F
00800713
F6E794E3
03000593
F59FF06F
03000593
00098513
000A00E7
FFF90913
FF2048E3
FFF40793
00045463
00000413
40878433
F49FF06F
00098513
000A00E7
F41FF06F
02000593
00098513
000A00E7
FFF40413
F49FF06F
00852703
00052783
00F77863
00452783
00E787B3
00B78023
00852783
00178793
00F52423
00008067
00452703
00052783
00170693
00D52223
00E787B3
00B78023
00008067
FA010113
05412423
01810793
00002A37
04912A23
05212823
05312623
05512223
05612023
03712E23
04112E23
04812C23
03812C23
00050493
00058913
00068B93
00F12A23
02500A93
02D00993
884A0A13
00500B13
00064583
00160413
02059A63
05C12083
05812403
05412483
05012903
04C12983
04812A03
04412A83
04012B03
03C12B83
03812C03
06010113
00008067
01558863
00048513
000900E7
1400006F
00414783
00012423
00010623
FF47F793
00F10223
00000713
00000693
00000613
03000593
02300513
00044783
00140413
00078863
05378E63
06B78063
06A78263
00060863
00414603
00866613
00C10223
00068863
00414683
0016E693
00D10223
00070863
00414703
00276713
00E10223
FD078713
0FF77713
00900693
06E6E063
00000613
00900593
00A00693
02C0006F
00100613
F95FF06F
00100693
F8DFF06F
00100713
F85FF06F
02D60633
00044783
00140413
00C70633
FD078713
0FF77513
FEA5F4E3
F9F78713
0FF77713
06EB6C63
FA978713
FCD70AE3
00C12423
02E00713
02E79463
00414783
00900693
0017E793
00F10223
00044783
00140413
FD078713
0FF77713
FEE6F8E3
07A00713
04E79663
00044783
00140413
00100713
07800693
00F6EE63
06200693
04F6EA63
1F578063
05800693
12D78A63
E80784E3
00040613
E75FF06F
FBF78713
0FF77713
F8EB66E3
FC978713
F81FF06F
06C00693
00000713
FAD79EE3
00044783
FAD796E3
00144783
00200713
00240413
FA5FF06F
F9D78613
0FF67613
01500693
FAC6EAE3
00261613
01460633
00062683
00068067
00A00793
00F12823
00200793
0EF71463
007B8693
FF86F693
0006A503
0046A583
00410613
00868B93
99DFF0EF
00410613
00090593
00048513
B95FF0EF
F65FF06F
00A00793
00F12823
00200793
04F71863
007B8B93
FF8BFB93
004BA583
000BA503
008B8C13
0005DC63
00A037B3
40B005B3
40F585B3
40A00533
01310623
00410613
945FF0EF
00410613
00090593
00048513
B3DFF0EF
000C0B93
F09FF06F
000BA503
004B8C13
00055663
40A00533
01310623
00410593
A8DFF0EF
FCDFF06F
00414703
00276713
00E10223
00000713
FA878793
0017B793
00279613
00414783
01000693
00D12823
FFB7F793
00C7E7B3
00F10223
F19FF06F
00100793
000BA503
00410593
004B8B93
00F71663
A39FF0EF
F21FF06F
A31FF0EF
F19FF06F
000BA503
00800793
00410593
00F12823
004B8C13
A15FF0EF
F55FF06F
000BC583
00048513
004B8C13
000900E7
F51FF06F
000BA783
00410613
00090593
00048513
00F12A23
A71FF0EF
01810793
004B8C13
00F12A23
F29FF06F
02500593
CE5FF06F
800007B7
20B7A223
800007B7
20A7A023
00008067
FC010113
02F12A23
800007B7
02B12223
2047A583
800007B7
02C12423
00050613
2007A503
02D12623
02410693
00112E23
02E12823
03012C23
03112E23
00D12623
BF9FF0EF
01C12083
04010113
00008067
04058C63
FE010113
FFF58593
00B12223
00A12423
5C400593
00410513
00112E23
00012623
BC5FF0EF
00C12683
00412703
00812783
00E6FE63
00D787B3
00078023
01C12083
00C12503
02010113
00008067
00E787B3
FE9FF06F
00000513
00008067
FC010113
02D12623
02C10693
00112E23
02E12823
02F12A23
03012C23
03112E23
00D12623
F7DFF0EF
01C12083
04010113
00008067
FE010113
00060693
00058613
00A12423
5EC00593
00810513
00112E23
00012623
B35FF0EF
00812783
00C12703
00E787B3
00078023
01C12083
00C12503
02010113
00008067
FC010113
02C12423
02810613
00112E23
02D12623
02E12823
02F12A23
03012C23
03112E23
00C12623
F95FF0EF
01C12083
04010113
00008067
FD010113
02812423
01712623
02112623
02912223
03212023
01312E23
01412C23
01512A23
01612823
01812423
01912223
00050B93
00058413
38069C63
000024B7
00060913
00050A13
8DC48493
12C5F863
000107B7
00058C13
10F67863
0FF00713
00C73733
00371713
00E657B3
00F484B3
0004C683
00E68733
02000693
40E687B3
00E68C63
00F41433
00EBD733
00F61933
00876C33
00FB9A33
01095B13
000B0593
000C0513
299000EF
00050493
000B0593
01091A93
000C0513
23D000EF
010ADA93
00050413
00050593
000A8513
1FD000EF
01049493
010A5713
00E4E733
00040993
00A77E63
01270733
FFF40993
01276863
00A77663
FFE40993
01270733
40A70433
000B0593
00040513
235000EF
00050493
000B0593
00040513
1DD000EF
010A1A13
00050413
00050593
01049493
000A8513
010A5A13
195000EF
0144EA33
00040613
00AA7C63
01490A33
FFF40613
012A6663
00AA7463
FFE40613
01099793
00C7E7B3
00000493
1300006F
010007B7
01000713
EEF66CE3
01800713
EF1FF06F
00068993
00061A63
00000593
00100513
169000EF
00050913
000107B7
12F97C63
0FF00793
0127F463
00800993
013957B3
00F484B3
0004C783
02000693
013787B3
40F68733
12F69263
41240433
00100493
01095A93
000A8593
00040513
165000EF
00050993
000A8593
00040513
01091B13
109000EF
010B5B13
00050413
00050593
000B0513
0C9000EF
01099993
010A5713
00E9E733
00040B93
00A77E63
01270733
FFF40B93
01276863
00A77663
FFE40B93
01270733
40A70433
000A8593
00040513
101000EF
00050993
000A8593
00040513
0A9000EF
010A1A13
00050413
00050593
01099993
000B0513
010A5A13
061000EF
0149EA33
00040613
00AA7C63
01490A33
FFF40613
012A6663
00AA7463
FFE40613
010B9793
00C7E7B3
00078513
00048593
02C12083
02812403
02412483
02012903
01C12983
01812A03
01412A83
01012B03
00C12B83
00812C03
00412C83
03010113
00008067
010007B7
01000993
ECF968E3
01800993
EC9FF06F
00E91933
00F459B3
00FBD7B3
00E41433
0087EAB3
01095413
00040593
00098513
00EB9A33
035000EF
00050493
00040593
00098513
01091B13
7D8000EF
010B5B13
00050993
00050593
000B0513
798000EF
01049493
010AD793
00F4E7B3
00098B93
00A7FE63
012787B3
FFF98B93
0127E863
00A7F663
FFE98B93
012787B3
40A789B3
00040593
00098513
7D0000EF
00040593
00050493
00098513
778000EF
010A9413
00050993
00050593
01049493
000B0513
01045413
730000EF
0084E433
00098793
00A47E63
01240433
FFF98793
01246863
00A47663
FFE98793
01240433
010B9493
40A40433
00F4E4B3
E01FF06F
1ED5EE63
000107B7
04F6F463
0FF00A93
00DAB733
00371713
000027B7
00E6D5B3
8DC78793
00B787B3
0007CA83
02000793
00EA8AB3
415784B3
03579663
00100793
E886E2E3
00CBB633
00164793
E79FF06F
010007B7
01000713
FCF6E0E3
01800713
FB9FF06F
01565CB3
009696B3
00DCECB3
015459B3
00941433
015BDAB3
008AEAB3
010CD413
00040593
00098513
00961933
6DC000EF
00050A13
00040593
00098513
010C9B13
680000EF
010B5B13
00050993
00050593
000B0513
640000EF
010A1A13
010AD713
00EA6733
00098C13
00A77E63
01970733
FFF98C13
01976863
00A77663
FFE98C13
01970733
40A709B3
00040593
00098513
678000EF
00040593
00050A13
00098513
620000EF
010A9413
00050993
00050593
010A1A13
000B0513
01045413
5D8000EF
008A6433
00098613
00A47E63
01940433
FFF98613
01946863
00A47663
FFE98613
01940433
010C1793
00010E37
00C7E7B3
FFFE0313
0067F8B3
00697333
40A40433
0107DE93
01095913
00088513
00030593
584000EF
00050813
00090593
00088513
574000EF
00050893
00030593
000E8513
564000EF
00050313
00090593
000E8513
554000EF
01085713
006888B3
01170733
00050693
00677463
01C506B3
01075513
00D506B3
02D46663
BCD412E3
00010537
FFF50513
00A77733
01071713
00A87833
009B9BB3
01070733
00000493
CCEBFAE3
FFF78793
B99FF06F
00000493
00000793
CC1FF06F
FD010113
02812423
02912223
03212023
01612823
02112623
01312E23
01412C23
01512A23
01712623
01812423
01912223
01A12023
00050913
00058B13
00050413
00058493
26069C63
00002AB7
00060A13
00068993
8DCA8A93
14C5F263
000107B7
12F67463
0FF00793
00C7F463
00800993
013657B3
00FA8AB3
000AC783
02000713
013787B3
40F709B3
00F70C63
013B15B3
00F957B3
01361A33
00B7E4B3
01391433
010A5A93
000A8593
00048513
4B8000EF
00050913
000A8593
010A1B13
00048513
45C000EF
010B5B13
00050593
000B0513
420000EF
01091913
01045793
00F967B3
00A7FA63
014787B3
0147E663
00A7F463
014787B3
40A784B3
000A8593
00048513
464000EF
00050913
000A8593
00048513
40C000EF
01041413
00050593
01091913
000B0513
01045413
3C8000EF
00896433
00A47A63
01440433
01446663
00A47463
01440433
40A40433
01345533
00000593
02C12083
02812403
02412483
02012903
01C12983
01812A03
01412A83
01012B03
00C12B83
00812C03
00412C83
00012D03
03010113
00008067
010007B7
01000993
EEF660E3
01800993
ED9FF06F
00061A63
00000593
00100513
374000EF
00050A13
000107B7
0EFA7A63
0FF00793
0147F463
00800993
013A57B3
00FA8AB3
000AC783
02000713
414B04B3
013787B3
40F709B3
ECF700E3
013A1A33
00FB5AB3
013B15B3
00F957B3
010A5493
00B7EB33
000A8513
00048593
360000EF
00048593
01391433
010A1B93
00050913
000A8513
300000EF
010BDB93
00050593
000B8513
2C4000EF
01091913
010B5793
00F967B3
00A7FA63
014787B3
0147E663
00A7F463
014787B3
40A78AB3
00048593
000A8513
308000EF
00050913
00048593
000A8513
2B0000EF
00050593
000B8513
278000EF
010B1593
01091913
0105D593
00B965B3
00A5FA63
014585B3
0145E663
00A5F463
014585B3
40A584B3
DFDFF06F
010007B7
01000993
F0FA6AE3
01800993
F0DFF06F
E8D5EAE3
000107B7
04F6FC63
0FF00A93
00DAB533
00351513
000027B7
00A6D733
8DC78793
00E787B3
0007CA83
02000793
00AA8AB3
41578A33
03579E63
0166E463
00C96A63
40C90433
40DB05B3
00893533
40A584B3
00040513
00048593
E39FF06F
010007B7
01000513
FAF6E8E3
01800513
FA9FF06F
014696B3
015657B3
00D7EC33
015B5D33
014B15B3
015954B3
010C5B13
00B4E4B3
000D0513
000B0593
01461CB3
208000EF
00050993
000B0593
000D0513
010C1B93
1AC000EF
010BDB93
00050593
01491433
00050913
000B8513
168000EF
01099993
0104D713
00E9E733
00090D13
00A77E63
01870733
FFF90D13
01876863
00A77663
FFE90D13
01870733
40A70933
000B0593
00090513
1A0000EF
00050993
000B0593
00090513
148000EF
00050913
00050593
000B8513
10C000EF
01049713
01099993
01075713
00E9E733
00090793
00A77E63
01870733
FFF90793
01876863
00A77663
FFE90793
01870733
00010EB7
010D1D13
00FD6D33
FFFE8793
00FD78B3
00FCF7B3
40A70733
010D5D13
010CDE13
00088513
00078593
0AC000EF
00050813
000E0593
00088513
09C000EF
00050893
00078593
000D0513
08C000EF
00050313
000E0593
000D0513
07C000EF
01085793
006888B3
011787B3
0067F463
01D50533
0107D593
00A585B3
00010537
FFF50513
00A7F7B3
01079793
00A87533
00A78533
00B76663
00B71E63
00A47C63
41950633
00C537B3
018787B3
40F585B3
00060513
40A40533
00A43433
40B705B3
408585B3
01559433
01455533
00A46533
0145D5B3
C65FF06F
00050613
00000513
0015F693
00068463
00C50533
0015D593
00161613
FE0596E3
00008067
06054063
0605C663
00058613
00050593
FFF00513
02060C63
00100693
00B67A63
00C05863
00161613
00169693
FEB66AE3
00000513
00C5E663
40C585B3
00D56533
0016D693
00165613
FE0696E3
00008067
00008293
FB5FF0EF
00058513
00028067
40A00533
00B04863
40B005B3
F9DFF06F
40B005B3
00008293
F91FF0EF
40A00533
00028067
00008293
0005CA63
00054C63
F79FF0EF
00058513
00028067
40B005B3
FE0558E3
40A00533
F61FF0EF
40B00533
00028067
FB010113
1EC00593
00000513
04112623
04912423
05212223
05312023
03412E23
03512C23
03612A23
03712823
03812623
ABCFF0EF
900007B7
03D00713
00002537
00E78023
84850993
84850513
AB4FF0EF
01498513
00010593
AA8FF0EF
910007B7
00600713
61616A37
00E78023
00000A93
161A0A13
00002BB7
90000937
000024B7
03098993
91000B37
00100C13
00010593
868B8513
01412023
01412223
A64FF0EF
00014783
00010593
868B8513
00178793
00F10023
00114783
001A8A93
00278793
00F100A3
00214783
00378793
00F10123
00314783
00478793
00F101A3
A24FF0EF
00094583
87048513
0FF5F593
A14FF0EF
00194583
87048513
0FF5F593
A04FF0EF
00294583
87048513
0FF5F593
9F4FF0EF
00394583
87048513
0FF5F593
9E4FF0EF
00494583
87048513
0FF5F593
9D4FF0EF
00594583
87048513
0FF5F593
9C4FF0EF
00694583
87048513
0FF5F593
9B4FF0EF
000A8593
00098513
9A8FF0EF
0C800513
018B0023
969FE0EF
0C800513
000B0023
95DFE0EF
F19FF06F
49520A0D
562D4353
6F6F4220
676E6974
00000A0D
3D667562
0A0D7025
00000000
3D667562
000A7325
0A0D7825
00000000
6E756F43
25203A74
00000A64
00000978
00000884
000007E4
000007E4
000007E4
000007E4
00000884
000007E4
000007E4
000007E4
000007E4
000007E4
0000095C
00000900
000007E4
000007E4
0000098C
000007E4
00000844
000007E4
000007E4
00000910
02020100
03030303
04040404
04040404
05050505
05050505
05050505
05050505
06060606
06060606
06060606
06060606
06060606
06060606
06060606
06060606
07070707
07070707
07070707
07070707
07070707
07070707
07070707
07070707
07070707
07070707
07070707
07070707
07070707
07070707
07070707
07070707
08080808
08080808
08080808
08080808
08080808
08080808
08080808
08080808
08080808
08080808
08080808
08080808
08080808
08080808
08080808
08080808
08080808
08080808
08080808
08080808
08080808
08080808
08080808
08080808
08080808
08080808
08080808
08080808
08080808
08080808
08080808
08080808
00000010
00000000
00527A03
01017C01
00020D1B
00000048
00000018
FFFFF138
000005D8
300E4400
9702886C
89018109
93049203
95069405
98089607
030B990A
C10A0270
C944C844
D344D244
D544D444
D744D644
D944D844
44000E44
0000000B
0000004C
00000064
FFFFF6C4
000004F0
300E4400
89028870
96049203
93018108
95069405
98099707
9A0B990A
0120030C
C844C10A
D244C944
D444D344
D644D544
D844D744
DA44D944
44000E44
0000000B
00000000
	 
